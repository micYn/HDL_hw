module wrapper(
    output wire layer1_enable1, layer1_enable2, layer1_enable3,
    output wire signed [35:0] output_feature_map1_pixel_layer1, output_feature_map2_pixel_layer1, output_feature_map3_pixel_layer1, output_feature_map4_pixel_layer1,
    output wire layer2_enable1, layer2_enable2, layer2_enable3, layer2_enable4,
    output wire signed [35:0] output_feature_map1_pixel_layer2, output_feature_map2_pixel_layer2, output_feature_map3_pixel_layer2, output_feature_map4_pixel_layer2,
    input wire signed [8:0] channel1_layer1, channel2_layer1, channel3_layer1, channel4_layer1,
                            channel1_layer2, channel2_layer2, channel3_layer2, channel4_layer2,
    input wire signed [15:0] weight111, weight112, weight113, weight114, weight115, weight116, weight117, weight118, weight119,
                             weight121, weight122, weight123, weight124, weight125, weight126, weight127, weight128, weight129,
                             weight131, weight132, weight133, weight134, weight135, weight136, weight137, weight138, weight139, 
                             weight141, weight142, weight143, weight144, weight145, weight146, weight147, weight148, weight149,

                             weight211, weight212, weight213, weight214, weight215, weight216, weight217, weight218, weight219,
                             weight221, weight222, weight223, weight224, weight225, weight226, weight227, weight228, weight229,
                             weight231, weight232, weight233, weight234, weight235, weight236, weight237, weight238, weight239, 
                             weight241, weight242, weight243, weight244, weight245, weight246, weight247, weight248, weight249,

                             weight311, weight312, weight313, weight314, weight315, weight316, weight317, weight318, weight319,
                             weight321, weight322, weight323, weight324, weight325, weight326, weight327, weight328, weight329,
                             weight331, weight332, weight333, weight334, weight335, weight336, weight337, weight338, weight339, 
                             weight341, weight342, weight343, weight344, weight345, weight346, weight347, weight348, weight349,

                             weight411, weight412, weight413, weight414, weight415, weight416, weight417, weight418, weight419,
                             weight421, weight422, weight423, weight424, weight425, weight426, weight427, weight428, weight429,
                             weight431, weight432, weight433, weight434, weight435, weight436, weight437, weight438, weight439, 
                             weight441, weight442, weight443, weight444, weight445, weight446, weight447, weight448, weight449,
    input wire signed [15:0] bias1, bias2, bias3, bias4,
    input wire clk,
    input wire rst
);
conv_layer1 conv_layer1_ins(layer1_enable1, layer1_enable2, layer1_enable3, output_feature_map1_pixel_layer1, output_feature_map2_pixel_layer1, output_feature_map3_pixel_layer1, output_feature_map4_pixel_layer1,
                                
                            channel1_layer1, channel2_layer1, channel3_layer1,
                            
                            weight111, weight112, weight113, weight114, weight115, weight116, weight117, weight118, weight119,
                            weight121, weight122, weight123, weight124, weight125, weight126, weight127, weight128, weight129,
                            weight131, weight132, weight133, weight134, weight135, weight136, weight137, weight138, weight139,

                            weight211, weight212, weight213, weight214, weight215, weight216, weight217, weight218, weight219,
                            weight221, weight222, weight223, weight224, weight225, weight226, weight227, weight228, weight229,
                            weight231, weight232, weight233, weight234, weight235, weight236, weight237, weight238, weight239,

                            weight311, weight312, weight313, weight314, weight315, weight316, weight317, weight318, weight319,
                            weight321, weight322, weight323, weight324, weight325, weight326, weight327, weight328, weight329,
                            weight331, weight332, weight333, weight334, weight335, weight336, weight337, weight338, weight339,

                            weight411, weight412, weight413, weight414, weight415, weight416, weight417, weight418, weight419,
                            weight421, weight422, weight423, weight424, weight425, weight426, weight427, weight428, weight429,
                            weight431, weight432, weight433, weight434, weight435, weight436, weight437, weight438, weight439,

                            bias1, bias2, bias3, bias4,

                            clk, rst);
    conv_layer2 conv_layer2_ins(layer2_enable1, layer2_enable2, layer2_enable3, layer2_enable4, output_feature_map1_pixel_layer2, output_feature_map2_pixel_layer2, output_feature_map3_pixel_layer2, output_feature_map4_pixel_layer2,
                                
                                channel1_layer2, channel2_layer2, channel3_layer2, channel4_layer2,
                                
                                weight111, weight112, weight113, weight114, weight115, weight116, weight117, weight118, weight119,
                                weight121, weight122, weight123, weight124, weight125, weight126, weight127, weight128, weight129,
                                weight131, weight132, weight133, weight134, weight135, weight136, weight137, weight138, weight139, 
                                weight141, weight142, weight143, weight144, weight145, weight146, weight147, weight148, weight149,

                                weight211, weight212, weight213, weight214, weight215, weight216, weight217, weight218, weight219,
                                weight221, weight222, weight223, weight224, weight225, weight226, weight227, weight228, weight229,
                                weight231, weight232, weight233, weight234, weight235, weight236, weight237, weight238, weight239, 
                                weight241, weight242, weight243, weight244, weight245, weight246, weight247, weight248, weight249,

                                weight311, weight312, weight313, weight314, weight315, weight316, weight317, weight318, weight319,
                                weight321, weight322, weight323, weight324, weight325, weight326, weight327, weight328, weight329,
                                weight331, weight332, weight333, weight334, weight335, weight336, weight337, weight338, weight339, 
                                weight341, weight342, weight343, weight344, weight345, weight346, weight347, weight348, weight349,

                                weight411, weight412, weight413, weight414, weight415, weight416, weight417, weight418, weight419,
                                weight421, weight422, weight423, weight424, weight425, weight426, weight427, weight428, weight429,
                                weight431, weight432, weight433, weight434, weight435, weight436, weight437, weight438, weight439, 
                                weight441, weight442, weight443, weight444, weight445, weight446, weight447, weight448, weight449,

                                bias1, bias2, bias3, bias4,

                                clk, rst);
endmodule